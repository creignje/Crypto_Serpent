LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Round IS
END ENTITY;

ARCHITECTURE Behavioral OF Round IS
BEGIN

END Behavioral;