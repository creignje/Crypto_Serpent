LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Linear_Transformation IS
END Linear_Transformation;

ARCHITECTURE Behavioral OF Linear_Transformation IS
BEGIN
END Behavioral;