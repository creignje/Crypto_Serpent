LIBRARY IEEE;

ENTITY Final_Permutation IS
END Final_Permutation;

ARCHITECTURE Behavioral OF Final_Permutation IS
BEGIN
END Behavioral;