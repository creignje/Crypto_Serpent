LIBRARY IEEE;

ENTITY tb_Final_Permutation IS
END tb_Final_Permutation;

ARCHITECTURE Behavioral OF tb_Final_Permutation IS
BEGIN
END Behavioral;