LIBRARY IEEE;

ENTITY tb_Initial_Permutation IS
END tb_Initial_Permutation;

ARCHITECTURE Behavioral OF tb_Initial_Permutation IS
BEGIN
END Behavioral;