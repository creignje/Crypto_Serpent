LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY tb_Linear_Transformation IS
END tb_Linear_Transformation;

ARCHITECTURE Behavioral OF tb_Linear_Transformation IS
BEGIN
END Behavioral;
