LIBRARY IEEE;

ENTITY Initial_Permutation IS
END Initial_Permutation;

ARCHITECTURE Behavioral OF Initial_Permutation IS
BEGIN
END Behavioral;