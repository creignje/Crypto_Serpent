LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Sbox0 IS
END Sbox0;

ARCHITECTURE Behavioral OF Sbox0 IS
BEGIN
END Behavioral;